//这是CostasLoop.v文件的程序清单
module Polar (
	rst,clk,din,
	di,dq,df); 
	
	input		rst;   //复位信号，高电平有效
	input		clk;   //FPGA系统时钟：8MHz
	input	 signed [7:0]	din;    //输入数据：8MHz
	output signed [25:0]	di;     //同步后的输出信号(同相支路)
	output signed [25:0]	dq;     //同步后的输出信号(正交支路)
	output signed [25:0]	df;     //环路滤波器输出数据
	
	//实例化NCO核所需的接口信号
	wire reset_n,out_valid,clken;
	wire [29:0] carrier;
	wire signed [9:0] sin,cos ;
	wire signed [29:0] frequency_df;
	wire signed [25:0] Loopout;
	assign reset_n = !rst;
	assign clken = 1'b1;
	//assign carrier=30'd268435456;//2MHz
	assign carrier=30'd53687091;//13421773;//100khz//268460000;//2.0002MHz
	
	assign frequency_df={{4{Loopout[25]}},Loopout};//根据NCO核接口，扩展为30位
	
	//实例化NCO核
   //Quartus提供的NCO核输出数据最小位宽为10比特，根据环路设计需求，只取高8比特参与后续运算	
	nco2m	u0 (
		.phi_inc_i (carrier),
		.clk (clk),
		.reset_n (reset_n),
		.clken (clken),
		.freq_mod_i (frequency_df),
		.fsin_o (sin),
		.fcos_o (cos),
		.out_valid (out_valid));
	
   //实例化NCO同相支路乘法运算器核
	wire signed [15:0] zi;	
   mult8_8 u1 (
	   .clock (clk),
		.dataa (sin[9:2]),
		.datab (din),
		.result (zi));
		
   //实例化NCO正交支路乘法运算器核	
	wire signed [15:0] zq;	
   mult8_8 u2 (
	   .clock (clk),
		.dataa (cos[9:2]),
		.datab (din),
		.result (zq));
		

   //实例化鉴相器同相支路低通滤波器核
	wire ast_sink_valid,ast_source_ready;
	wire [1:0] ast_source_error;
	wire [1:0] ast_sink_error;
	assign ast_sink_valid=1'b1;
	assign ast_source_ready=1'b1;
	assign ast_sink_error=2'd0;
	wire sink_readyi,source_validi;
	wire [1:0] source_errori;
	wire signed [26:0] yi;	
   fir_lpf u3(
		.clk (clk),
		.reset_n (reset_n),
		.ast_sink_data (zi[14:0]),
		.ast_sink_valid (ast_sink_valid),
		.ast_source_ready (ast_source_ready),
		.ast_sink_error (ast_sink_error),
		.ast_source_data (yi),
		.ast_sink_ready (sink_readyi),
		.ast_source_valid (source_validi),
		.ast_source_error (source_errori));


   //实例化鉴相器正交支路低通滤波器核
	wire sink_readyq,source_validq;
	wire [1:0] source_errorq;
	wire signed [26:0] yq;	
   fir_lpf u4(
		.clk (clk),
		.reset_n (reset_n),
		.ast_sink_data (zq[14:0]),
		.ast_sink_valid (ast_sink_valid),
		.ast_source_ready (ast_source_ready),
		.ast_sink_error (ast_sink_error),
		.ast_source_data (yq),
		.ast_sink_ready (sink_readyq),
		.ast_source_valid (source_validq),
		.ast_source_error (source_erroriq));
		
		
   //根据同相支路的符号位，取正交支路数据（或取反）作为鉴相器输出
	reg signed [26:0] pd;
	always @(posedge clk or posedge rst)
		if (rst)
		   pd <= 0;
		else
			if	(yi[26]==1'b1)
				pd <= -yq;
			else
				pd <= yq;
			
	//实例化环路滤波器模块	
   LoopFilter u5(
	   .rst (rst),
		.clk (clk),
		.pd  (pd[26:1]),
		.frequency_df(Loopout));
		
	//将环路滤波器数据送至输出端口查看	
	assign df = Loopout;
	assign di = yi[26:1];
	assign dq = yq[26:1];
	
endmodule
